module bridgetop(HCLK,HRESET,PENABLE,PWRITE,PSEL,PADDR,PWDATA,HREADYOUT,HWRITE,HREADYIN,HWDATA,HADDR,HTRANS);

input HCLK,HRESET,HWRITE,HREADYIN;
input[1:0] HTRANS;
input[31:0] HWDATA,HADDR;

output wire PENABLE,PWRITE,HREADYOUT;
output wire [2:0] PSEL;
output wire [31:0] PADDR,PWDATA;

wire w1,w7;
wire[2:0]w2;
wire[31:0]w3,w4,w5,w6;

ahbslave ahb(.HCLK(HCLK),.HWRITE(HWRITE),.HRESET(HRESET),.HREADYIN(HREADYIN),.HTRANS(HTRANS),.HWDATA(HWDATA),.HADDR(HADDR),.VALID(w1),.TEMP_SEL(w2),.PIPEA0(w3),.PIPEA1(w4),.PIPED0(w5),.PIPED1(w6), .HWRITEREG(w7));

fsmcontroller fsm(.HCLK(HCLK),.HRESETn(HRESET),.VALID(w1),.HWDATA0(w5),.HWDATA1(w6),.HADDR0(w3),.HADDR1(w4),.TEMP(w2),.PENABLE(PENABLE),.PWRITE(PWRITE),.HREADOUT(HREADYOUT),.PSEL(PSEL),.PADDR(PADDR),.PWDATA(PWDATA),.HWRITE(HWRITE),.HWRITEREG(w7));


endmodule
